module csr(
    input logic clk,
    input logic rst_n,
    // 现在先不写了x
);

endmodule